BLUE
0 0 0 0 0 r h 
0 0 0 0 0 r h 
0 0 0 0 0 r h 
0 0 0 0 0 r h 
336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 336 0 
0